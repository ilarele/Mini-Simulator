*7 9
V 1 0 PULSE(4 12 5 2 3 5 19)
R 1 2 1
R 2 3 2
R 3 4 3
R 4 5 4
R 5 6 5
R 0 6 6
R 5 2 7
R 6 4 8
.TRAN 0.2 40
.PLOT TRAN V(4,2)
