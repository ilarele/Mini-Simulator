*3 3
V 1 0 PULSE(3 10 2 2 2 3 10)
C 1 2 3
R 2 0 1
.TRAN 0.2 40
.PLOT TRAN V(1,2)
