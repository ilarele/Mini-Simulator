*4 5
V 1 0 PULSE(3 10 1 3 5 5 20)
C 2 0 3
C 2 3 3
R 1 2 5
R 0 3 1
.TRAN 0.2 40
.PLOT TRAN V(1,3)