*5 6
V 1 0 PULSE(5 10 0 2 1 5 10)
R 1 2 2
C 2 3 10
R 3 4 10
R 1 4 2
C 0 4 10
.TRAN 0.2 40
.PLOT TRAN V(3,4)